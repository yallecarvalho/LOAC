{"devices":{"dev0":{"label":"J1","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J1","order":0,"position":{"x":12,"y":12}},"dev1":{"label":"J2","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J2","order":1,"position":{"x":12,"y":62}},"dev2":{"label":"J3","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J3","order":2,"position":{"x":12,"y":112}},"dev3":{"label":"J4","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J4","order":3,"position":{"x":12,"y":162}},"dev4":{"label":"J5","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J5","order":4,"position":{"x":12,"y":212}},"dev5":{"label":"J6","type":"Button","propagation":0,"numbase":"hex","bits":1,"net":"J6","order":5,"position":{"x":12,"y":262}},"dev6":{"label":"saida_alarme","type":"Lamp","propagation":0,"numbase":"hex","bits":1,"net":"saida_alarme","order":6,"position":{"x":422,"y":120}},"dev11":{"label":"$or$alarme.sv:5$6","type":"Or","propagation":1,"source_positions":[{"name":"alarme.sv","from":{"line":5,"column":32},"to":{"line":5,"column":59}}],"bits":1,"inputs":6,"position":{"x":142,"y":87}}},"connectors":[{"from":{"id":"dev11","port":"out"},"to":{"id":"dev6","port":"in"},"name":"saida_alarme"},{"from":{"id":"dev5","port":"out"},"to":{"id":"dev11","port":"in6"},"name":"J6","vertices":[{"x":92,"y":277},{"x":102,"y":267},{"x":102,"y":185}]},{"from":{"id":"dev4","port":"out"},"to":{"id":"dev11","port":"in5"},"name":"J5","vertices":[{"x":92,"y":217},{"x":92,"y":169}]},{"from":{"id":"dev3","port":"out"},"to":{"id":"dev11","port":"in4"},"name":"J4","vertices":[{"x":82,"y":167},{"x":82,"y":153},{"x":92,"y":143}]},{"from":{"id":"dev2","port":"out"},"to":{"id":"dev11","port":"in3"},"name":"J3"},{"from":{"id":"dev0","port":"out"},"to":{"id":"dev11","port":"in1"},"name":"J1","vertices":[{"x":92,"y":37},{"x":92,"y":85}]},{"from":{"id":"dev1","port":"out"},"to":{"id":"dev11","port":"in2"},"name":"J2","vertices":[{"x":82,"y":87},{"x":82,"y":101},{"x":92,"y":111}]}],"subcircuits":{}}